module SDRAM_Ctrl(

);


endmodule