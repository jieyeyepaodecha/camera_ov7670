module FIFO_Write(
input	wire	sclk,
input	wire	rst_n,
input	wire	[15:0]  FIFO_in_data
);


endmodule