module FIFO_Write(
input	wire	sclk,
input	wire	rst_n
);


endmodule