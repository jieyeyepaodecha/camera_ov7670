module FIFO_Read(
input	wire	sclk,
input	wire	rst_n,
input	wire	[15:0]  FIFO_Data,
output	reg		FIFO_Read_en
);


endmodule